// nios_cpu.v

// Generated using ACDS version 16.1 200

`timescale 1 ps / 1 ps
module nios_cpu (
		input  wire        clk_clk,                                //                  clk.clk
		input  wire        dac_spi1_MISO,                          //             dac_spi1.MISO
		output wire        dac_spi1_MOSI,                          //                     .MOSI
		output wire        dac_spi1_SCLK,                          //                     .SCLK
		output wire        dac_spi1_SS_n,                          //                     .SS_n
		input  wire [31:0] exfifo_if_d_export,                     //          exfifo_if_d.export
		output wire        exfifo_if_rd_export,                    //         exfifo_if_rd.export
		input  wire        exfifo_if_rdempty_export,               //    exfifo_if_rdempty.export
		output wire [31:0] exfifo_of_d_export,                     //          exfifo_of_d.export
		output wire        exfifo_of_wr_export,                    //         exfifo_of_wr.export
		input  wire        exfifo_of_wrfull_export,                //     exfifo_of_wrfull.export
		output wire        exfifo_rst_export,                      //           exfifo_rst.export
		input  wire        fpga_spi0_MISO,                         //            fpga_spi0.MISO
		output wire        fpga_spi0_MOSI,                         //                     .MOSI
		output wire        fpga_spi0_SCLK,                         //                     .SCLK
		output wire [7:0]  fpga_spi0_SS_n,                         //                     .SS_n
		input  wire [7:0]  gpi0_export,                            //                 gpi0.export
		output wire [7:0]  gpio0_export,                           //                gpio0.export
		input  wire [63:0] pll_recfg_from_pll_0_reconfig_from_pll, // pll_recfg_from_pll_0.reconfig_from_pll
		input  wire [63:0] pll_recfg_from_pll_1_reconfig_from_pll, // pll_recfg_from_pll_1.reconfig_from_pll
		input  wire [63:0] pll_recfg_from_pll_2_reconfig_from_pll, // pll_recfg_from_pll_2.reconfig_from_pll
		input  wire [63:0] pll_recfg_from_pll_3_reconfig_from_pll, // pll_recfg_from_pll_3.reconfig_from_pll
		input  wire [63:0] pll_recfg_from_pll_4_reconfig_from_pll, // pll_recfg_from_pll_4.reconfig_from_pll
		input  wire [63:0] pll_recfg_from_pll_5_reconfig_from_pll, // pll_recfg_from_pll_5.reconfig_from_pll
		output wire [63:0] pll_recfg_to_pll_0_reconfig_to_pll,     //   pll_recfg_to_pll_0.reconfig_to_pll
		output wire [63:0] pll_recfg_to_pll_1_reconfig_to_pll,     //   pll_recfg_to_pll_1.reconfig_to_pll
		output wire [63:0] pll_recfg_to_pll_2_reconfig_to_pll,     //   pll_recfg_to_pll_2.reconfig_to_pll
		output wire [63:0] pll_recfg_to_pll_3_reconfig_to_pll,     //   pll_recfg_to_pll_3.reconfig_to_pll
		output wire [63:0] pll_recfg_to_pll_4_reconfig_to_pll,     //   pll_recfg_to_pll_4.reconfig_to_pll
		output wire [63:0] pll_recfg_to_pll_5_reconfig_to_pll,     //   pll_recfg_to_pll_5.reconfig_to_pll
		output wire [31:0] pll_rst_export,                         //              pll_rst.export
		input  wire [3:0]  pllcfg_cmd_export,                      //           pllcfg_cmd.export
		input  wire        pllcfg_spi_MISO,                        //           pllcfg_spi.MISO
		output wire        pllcfg_spi_MOSI,                        //                     .MOSI
		output wire        pllcfg_spi_SCLK,                        //                     .SCLK
		output wire        pllcfg_spi_SS_n,                        //                     .SS_n
		output wire [9:0]  pllcfg_stat_export,                     //          pllcfg_stat.export
		inout  wire        scl_export,                             //                  scl.export
		inout  wire        sda_export                              //                  sda.export
	);

	wire         nios2_cpu_debug_reset_request_reset;                            // nios2_cpu:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire  [31:0] nios2_cpu_data_master_readdata;                                 // mm_interconnect_0:nios2_cpu_data_master_readdata -> nios2_cpu:d_readdata
	wire         nios2_cpu_data_master_waitrequest;                              // mm_interconnect_0:nios2_cpu_data_master_waitrequest -> nios2_cpu:d_waitrequest
	wire         nios2_cpu_data_master_debugaccess;                              // nios2_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_cpu_data_master_debugaccess
	wire  [16:0] nios2_cpu_data_master_address;                                  // nios2_cpu:d_address -> mm_interconnect_0:nios2_cpu_data_master_address
	wire   [3:0] nios2_cpu_data_master_byteenable;                               // nios2_cpu:d_byteenable -> mm_interconnect_0:nios2_cpu_data_master_byteenable
	wire         nios2_cpu_data_master_read;                                     // nios2_cpu:d_read -> mm_interconnect_0:nios2_cpu_data_master_read
	wire         nios2_cpu_data_master_write;                                    // nios2_cpu:d_write -> mm_interconnect_0:nios2_cpu_data_master_write
	wire  [31:0] nios2_cpu_data_master_writedata;                                // nios2_cpu:d_writedata -> mm_interconnect_0:nios2_cpu_data_master_writedata
	wire  [31:0] nios2_cpu_instruction_master_readdata;                          // mm_interconnect_0:nios2_cpu_instruction_master_readdata -> nios2_cpu:i_readdata
	wire         nios2_cpu_instruction_master_waitrequest;                       // mm_interconnect_0:nios2_cpu_instruction_master_waitrequest -> nios2_cpu:i_waitrequest
	wire  [16:0] nios2_cpu_instruction_master_address;                           // nios2_cpu:i_address -> mm_interconnect_0:nios2_cpu_instruction_master_address
	wire         nios2_cpu_instruction_master_read;                              // nios2_cpu:i_read -> mm_interconnect_0:nios2_cpu_instruction_master_read
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;       // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;    // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect;      // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_chipselect -> Av_FIFO_Int_0:chipselect
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata;        // Av_FIFO_Int_0:readdata -> mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_readdata
	wire   [1:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address;         // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_address -> Av_FIFO_Int_0:address
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read;            // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_read -> Av_FIFO_Int_0:read
	wire         mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write;           // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_write -> Av_FIFO_Int_0:write
	wire  [31:0] mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata;       // mm_interconnect_0:Av_FIFO_Int_0_avalon_slave_0_writedata -> Av_FIFO_Int_0:writedata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect;    // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_chipselect -> i2c_opencores_0:wb_stb_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata;      // i2c_opencores_0:wb_dat_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest;   // i2c_opencores_0:wb_ack_o -> mm_interconnect_0:i2c_opencores_0_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address;       // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_address -> i2c_opencores_0:wb_adr_i
	wire         mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write;         // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_write -> i2c_opencores_0:wb_we_i
	wire   [7:0] mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata;     // mm_interconnect_0:i2c_opencores_0_avalon_slave_0_writedata -> i2c_opencores_0:wb_dat_i
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;          // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;           // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata;           // nios2_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios2_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest;        // nios2_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess;        // mm_interconnect_0:nios2_cpu_debug_mem_slave_debugaccess -> nios2_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_address;            // mm_interconnect_0:nios2_cpu_debug_mem_slave_address -> nios2_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_read;               // mm_interconnect_0:nios2_cpu_debug_mem_slave_read -> nios2_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable;         // mm_interconnect_0:nios2_cpu_debug_mem_slave_byteenable -> nios2_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_cpu_debug_mem_slave_write;              // mm_interconnect_0:nios2_cpu_debug_mem_slave_write -> nios2_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata;          // mm_interconnect_0:nios2_cpu_debug_mem_slave_writedata -> nios2_cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata;    // pll_reconfig_0:mgmt_readdata -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest; // pll_reconfig_0:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_address -> pll_reconfig_0:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_read -> pll_reconfig_0:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_write -> pll_reconfig_0:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_0_mgmt_avalon_slave_writedata -> pll_reconfig_0:mgmt_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata;    // pll_reconfig_5:mgmt_readdata -> mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest; // pll_reconfig_5:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_address -> pll_reconfig_5:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_read -> pll_reconfig_5:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_write -> pll_reconfig_5:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_5_mgmt_avalon_slave_writedata -> pll_reconfig_5:mgmt_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata;    // pll_reconfig_4:mgmt_readdata -> mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest; // pll_reconfig_4:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_address -> pll_reconfig_4:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_read -> pll_reconfig_4:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_write -> pll_reconfig_4:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_4_mgmt_avalon_slave_writedata -> pll_reconfig_4:mgmt_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata;    // pll_reconfig_3:mgmt_readdata -> mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest; // pll_reconfig_3:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_address -> pll_reconfig_3:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_read -> pll_reconfig_3:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_write -> pll_reconfig_3:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_3_mgmt_avalon_slave_writedata -> pll_reconfig_3:mgmt_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata;    // pll_reconfig_2:mgmt_readdata -> mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest; // pll_reconfig_2:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_address -> pll_reconfig_2:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_read -> pll_reconfig_2:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_write -> pll_reconfig_2:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_2_mgmt_avalon_slave_writedata -> pll_reconfig_2:mgmt_writedata
	wire  [31:0] mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata;    // pll_reconfig_1:mgmt_readdata -> mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_readdata
	wire         mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest; // pll_reconfig_1:mgmt_waitrequest -> mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_waitrequest
	wire   [5:0] mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address;     // mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_address -> pll_reconfig_1:mgmt_address
	wire         mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read;        // mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_read -> pll_reconfig_1:mgmt_read
	wire         mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write;       // mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_write -> pll_reconfig_1:mgmt_write
	wire  [31:0] mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata;   // mm_interconnect_0:pll_reconfig_1_mgmt_avalon_slave_writedata -> pll_reconfig_1:mgmt_writedata
	wire         mm_interconnect_0_oc_mem_s1_chipselect;                         // mm_interconnect_0:oc_mem_s1_chipselect -> oc_mem:chipselect
	wire  [31:0] mm_interconnect_0_oc_mem_s1_readdata;                           // oc_mem:readdata -> mm_interconnect_0:oc_mem_s1_readdata
	wire  [12:0] mm_interconnect_0_oc_mem_s1_address;                            // mm_interconnect_0:oc_mem_s1_address -> oc_mem:address
	wire   [3:0] mm_interconnect_0_oc_mem_s1_byteenable;                         // mm_interconnect_0:oc_mem_s1_byteenable -> oc_mem:byteenable
	wire         mm_interconnect_0_oc_mem_s1_write;                              // mm_interconnect_0:oc_mem_s1_write -> oc_mem:write
	wire  [31:0] mm_interconnect_0_oc_mem_s1_writedata;                          // mm_interconnect_0:oc_mem_s1_writedata -> oc_mem:writedata
	wire         mm_interconnect_0_oc_mem_s1_clken;                              // mm_interconnect_0:oc_mem_s1_clken -> oc_mem:clken
	wire         mm_interconnect_0_gpio_0_s1_chipselect;                         // mm_interconnect_0:gpio_0_s1_chipselect -> gpio_0:chipselect
	wire  [31:0] mm_interconnect_0_gpio_0_s1_readdata;                           // gpio_0:readdata -> mm_interconnect_0:gpio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_gpio_0_s1_address;                            // mm_interconnect_0:gpio_0_s1_address -> gpio_0:address
	wire         mm_interconnect_0_gpio_0_s1_write;                              // mm_interconnect_0:gpio_0_s1_write -> gpio_0:write_n
	wire  [31:0] mm_interconnect_0_gpio_0_s1_writedata;                          // mm_interconnect_0:gpio_0_s1_writedata -> gpio_0:writedata
	wire  [31:0] mm_interconnect_0_gpi_0_s1_readdata;                            // gpi_0:readdata -> mm_interconnect_0:gpi_0_s1_readdata
	wire   [1:0] mm_interconnect_0_gpi_0_s1_address;                             // mm_interconnect_0:gpi_0_s1_address -> gpi_0:address
	wire  [31:0] mm_interconnect_0_pllcfg_command_s1_readdata;                   // PLLCFG_Command:readdata -> mm_interconnect_0:PLLCFG_Command_s1_readdata
	wire   [1:0] mm_interconnect_0_pllcfg_command_s1_address;                    // mm_interconnect_0:PLLCFG_Command_s1_address -> PLLCFG_Command:address
	wire         mm_interconnect_0_pllcfg_status_s1_chipselect;                  // mm_interconnect_0:PLLCFG_Status_s1_chipselect -> PLLCFG_Status:chipselect
	wire  [31:0] mm_interconnect_0_pllcfg_status_s1_readdata;                    // PLLCFG_Status:readdata -> mm_interconnect_0:PLLCFG_Status_s1_readdata
	wire   [1:0] mm_interconnect_0_pllcfg_status_s1_address;                     // mm_interconnect_0:PLLCFG_Status_s1_address -> PLLCFG_Status:address
	wire         mm_interconnect_0_pllcfg_status_s1_write;                       // mm_interconnect_0:PLLCFG_Status_s1_write -> PLLCFG_Status:write_n
	wire  [31:0] mm_interconnect_0_pllcfg_status_s1_writedata;                   // mm_interconnect_0:PLLCFG_Status_s1_writedata -> PLLCFG_Status:writedata
	wire         mm_interconnect_0_pll_rst_s1_chipselect;                        // mm_interconnect_0:PLL_RST_s1_chipselect -> PLL_RST:chipselect
	wire  [31:0] mm_interconnect_0_pll_rst_s1_readdata;                          // PLL_RST:readdata -> mm_interconnect_0:PLL_RST_s1_readdata
	wire   [1:0] mm_interconnect_0_pll_rst_s1_address;                           // mm_interconnect_0:PLL_RST_s1_address -> PLL_RST:address
	wire         mm_interconnect_0_pll_rst_s1_write;                             // mm_interconnect_0:PLL_RST_s1_write -> PLL_RST:write_n
	wire  [31:0] mm_interconnect_0_pll_rst_s1_writedata;                         // mm_interconnect_0:PLL_RST_s1_writedata -> PLL_RST:writedata
	wire         mm_interconnect_0_fpga_spi0_spi_control_port_chipselect;        // mm_interconnect_0:fpga_spi0_spi_control_port_chipselect -> fpga_spi0:spi_select
	wire  [15:0] mm_interconnect_0_fpga_spi0_spi_control_port_readdata;          // fpga_spi0:data_to_cpu -> mm_interconnect_0:fpga_spi0_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_fpga_spi0_spi_control_port_address;           // mm_interconnect_0:fpga_spi0_spi_control_port_address -> fpga_spi0:mem_addr
	wire         mm_interconnect_0_fpga_spi0_spi_control_port_read;              // mm_interconnect_0:fpga_spi0_spi_control_port_read -> fpga_spi0:read_n
	wire         mm_interconnect_0_fpga_spi0_spi_control_port_write;             // mm_interconnect_0:fpga_spi0_spi_control_port_write -> fpga_spi0:write_n
	wire  [15:0] mm_interconnect_0_fpga_spi0_spi_control_port_writedata;         // mm_interconnect_0:fpga_spi0_spi_control_port_writedata -> fpga_spi0:data_from_cpu
	wire         mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect;       // mm_interconnect_0:PLLCFG_SPI_spi_control_port_chipselect -> PLLCFG_SPI:spi_select
	wire  [15:0] mm_interconnect_0_pllcfg_spi_spi_control_port_readdata;         // PLLCFG_SPI:data_to_cpu -> mm_interconnect_0:PLLCFG_SPI_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_pllcfg_spi_spi_control_port_address;          // mm_interconnect_0:PLLCFG_SPI_spi_control_port_address -> PLLCFG_SPI:mem_addr
	wire         mm_interconnect_0_pllcfg_spi_spi_control_port_read;             // mm_interconnect_0:PLLCFG_SPI_spi_control_port_read -> PLLCFG_SPI:read_n
	wire         mm_interconnect_0_pllcfg_spi_spi_control_port_write;            // mm_interconnect_0:PLLCFG_SPI_spi_control_port_write -> PLLCFG_SPI:write_n
	wire  [15:0] mm_interconnect_0_pllcfg_spi_spi_control_port_writedata;        // mm_interconnect_0:PLLCFG_SPI_spi_control_port_writedata -> PLLCFG_SPI:data_from_cpu
	wire         mm_interconnect_0_dac_spi1_spi_control_port_chipselect;         // mm_interconnect_0:dac_spi1_spi_control_port_chipselect -> dac_spi1:spi_select
	wire  [15:0] mm_interconnect_0_dac_spi1_spi_control_port_readdata;           // dac_spi1:data_to_cpu -> mm_interconnect_0:dac_spi1_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_dac_spi1_spi_control_port_address;            // mm_interconnect_0:dac_spi1_spi_control_port_address -> dac_spi1:mem_addr
	wire         mm_interconnect_0_dac_spi1_spi_control_port_read;               // mm_interconnect_0:dac_spi1_spi_control_port_read -> dac_spi1:read_n
	wire         mm_interconnect_0_dac_spi1_spi_control_port_write;              // mm_interconnect_0:dac_spi1_spi_control_port_write -> dac_spi1:write_n
	wire  [15:0] mm_interconnect_0_dac_spi1_spi_control_port_writedata;          // mm_interconnect_0:dac_spi1_spi_control_port_writedata -> dac_spi1:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                       // i2c_opencores_0:wb_inta_o -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                       // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                       // fpga_spi0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                       // PLLCFG_SPI:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                       // dac_spi1:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_cpu_irq_irq;                                              // irq_mapper:sender_irq -> nios2_cpu:irq
	wire         rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [Av_FIFO_Int_0:rsi_nrst, mm_interconnect_0:Av_FIFO_Int_0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [PLLCFG_Command:reset_n, PLLCFG_SPI:reset_n, PLLCFG_Status:reset_n, PLL_RST:reset_n, dac_spi1:reset_n, fpga_spi0:reset_n, gpi_0:reset_n, gpio_0:reset_n, i2c_opencores_0:wb_rst_i, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_cpu_reset_reset_bridge_in_reset_reset, nios2_cpu:reset_n, oc_mem:reset, pll_reconfig_0:mgmt_reset, pll_reconfig_1:mgmt_reset, pll_reconfig_2:mgmt_reset, pll_reconfig_3:mgmt_reset, pll_reconfig_4:mgmt_reset, pll_reconfig_5:mgmt_reset, rst_translator:in_reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                         // rst_controller_001:reset_req -> [nios2_cpu:reset_req, oc_mem:reset_req, rst_translator:reset_req_in]

	avfifo #(
		.width (32)
	) av_fifo_int_0 (
		.clk            (clk_clk),                                                   //          clock.clk
		.address        (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chipselect     (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect), //               .chipselect
		.write          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),      //               .write
		.writedata      (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),  //               .writedata
		.read           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),       //               .read
		.readdata       (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),   //               .readdata
		.rsi_nrst       (~rst_controller_reset_out_reset),                           //          reset.reset_n
		.coe_if_d       (exfifo_if_d_export),                                        //       cnd_if_d.export
		.coe_if_rd      (exfifo_if_rd_export),                                       //      cnd_if_rd.export
		.coe_of_wrfull  (exfifo_of_wrfull_export),                                   //  cnd_of_wrfull.export
		.coe_of_wr      (exfifo_of_wr_export),                                       //      cnd_of_wr.export
		.coe_of_d       (exfifo_of_d_export),                                        //       cnd_of_d.export
		.coe_if_rdempty (exfifo_if_rdempty_export),                                  // cnd_if_rdempty.export
		.coe_fifo_rst   (exfifo_rst_export)                                          //   cnd_fifo_rst.export
	);

	nios_cpu_PLLCFG_Command pllcfg_command (
		.clk      (clk_clk),                                      //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_pllcfg_command_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pllcfg_command_s1_readdata), //                    .readdata
		.in_port  (pllcfg_cmd_export)                             // external_connection.export
	);

	nios_cpu_PLLCFG_SPI pllcfg_spi (
		.clk           (clk_clk),                                                  //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                      //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_pllcfg_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_pllcfg_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_pllcfg_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_pllcfg_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_pllcfg_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver3_irq),                                 //              irq.irq
		.MISO          (pllcfg_spi_MISO),                                          //         external.export
		.MOSI          (pllcfg_spi_MOSI),                                          //                 .export
		.SCLK          (pllcfg_spi_SCLK),                                          //                 .export
		.SS_n          (pllcfg_spi_SS_n)                                           //                 .export
	);

	nios_cpu_PLLCFG_Status pllcfg_status (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pllcfg_status_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pllcfg_status_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pllcfg_status_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pllcfg_status_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pllcfg_status_s1_readdata),   //                    .readdata
		.out_port   (pllcfg_stat_export)                             // external_connection.export
	);

	nios_cpu_PLL_RST pll_rst (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_pll_rst_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pll_rst_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pll_rst_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pll_rst_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pll_rst_s1_readdata),   //                    .readdata
		.out_port   (pll_rst_export)                           // external_connection.export
	);

	nios_cpu_dac_spi1 dac_spi1 (
		.clk           (clk_clk),                                                //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                    //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_dac_spi1_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_dac_spi1_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_dac_spi1_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_dac_spi1_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_dac_spi1_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_dac_spi1_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver4_irq),                               //              irq.irq
		.MISO          (dac_spi1_MISO),                                          //         external.export
		.MOSI          (dac_spi1_MOSI),                                          //                 .export
		.SCLK          (dac_spi1_SCLK),                                          //                 .export
		.SS_n          (dac_spi1_SS_n)                                           //                 .export
	);

	nios_cpu_fpga_spi0 fpga_spi0 (
		.clk           (clk_clk),                                                 //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_fpga_spi0_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_fpga_spi0_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_fpga_spi0_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_fpga_spi0_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_fpga_spi0_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_fpga_spi0_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                //              irq.irq
		.MISO          (fpga_spi0_MISO),                                          //         external.export
		.MOSI          (fpga_spi0_MOSI),                                          //                 .export
		.SCLK          (fpga_spi0_SCLK),                                          //                 .export
		.SS_n          (fpga_spi0_SS_n)                                           //                 .export
	);

	nios_cpu_gpi_0 gpi_0 (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_gpi_0_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gpi_0_s1_readdata), //                    .readdata
		.in_port  (gpi0_export)                          // external_connection.export
	);

	nios_cpu_gpio_0 gpio_0 (
		.clk        (clk_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_gpio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpio_0_s1_readdata),   //                    .readdata
		.out_port   (gpio0_export)                            // external_connection.export
	);

	i2c_opencores i2c_opencores_0 (
		.wb_clk_i   (clk_clk),                                                      //            clock.clk
		.wb_rst_i   (rst_controller_001_reset_out_reset),                           //      clock_reset.reset
		.scl_pad_io (scl_export),                                                   //       export_scl.export
		.sda_pad_io (sda_export),                                                   //       export_sda.export
		.wb_adr_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_mapper_receiver0_irq)                                      // interrupt_sender.irq
	);

	nios_cpu_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	nios_cpu_nios2_cpu nios2_cpu (
		.clk                                 (clk_clk),                                                 //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios2_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios2_cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                         // custom_instruction_master.readra
	);

	nios_cpu_oc_mem oc_mem (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_oc_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_oc_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_oc_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_oc_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_oc_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_oc_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_oc_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_0 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_0_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_0_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_1 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_1_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_1_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_2 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_2_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_2_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_3 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_3_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_3_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_4 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_4_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_4_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	altera_pll_reconfig_top #(
		.device_family       ("Cyclone V"),
		.ENABLE_MIF          (0),
		.MIF_FILE_NAME       (""),
		.ENABLE_BYTEENABLE   (0),
		.BYTEENABLE_WIDTH    (4),
		.RECONFIG_ADDR_WIDTH (6),
		.RECONFIG_DATA_WIDTH (32),
		.reconf_width        (64),
		.WAIT_FOR_LOCK       (1)
	) pll_reconfig_5 (
		.mgmt_clk          (clk_clk),                                                        //          mgmt_clk.clk
		.mgmt_reset        (rst_controller_001_reset_out_reset),                             //        mgmt_reset.reset
		.mgmt_waitrequest  (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest), // mgmt_avalon_slave.waitrequest
		.mgmt_read         (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read),        //                  .read
		.mgmt_write        (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write),       //                  .write
		.mgmt_readdata     (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata),    //                  .readdata
		.mgmt_address      (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address),     //                  .address
		.mgmt_writedata    (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata),   //                  .writedata
		.reconfig_to_pll   (pll_recfg_to_pll_5_reconfig_to_pll),                             //   reconfig_to_pll.reconfig_to_pll
		.reconfig_from_pll (pll_recfg_from_pll_5_reconfig_from_pll),                         // reconfig_from_pll.reconfig_from_pll
		.mgmt_byteenable   (4'b0000)                                                         //       (terminated)
	);

	nios_cpu_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                   (clk_clk),                                                        //                                 clk_0_clk.clk
		.Av_FIFO_Int_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                 // Av_FIFO_Int_0_reset_reset_bridge_in_reset.reset
		.nios2_cpu_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                             //     nios2_cpu_reset_reset_bridge_in_reset.reset
		.nios2_cpu_data_master_address                   (nios2_cpu_data_master_address),                                  //                     nios2_cpu_data_master.address
		.nios2_cpu_data_master_waitrequest               (nios2_cpu_data_master_waitrequest),                              //                                          .waitrequest
		.nios2_cpu_data_master_byteenable                (nios2_cpu_data_master_byteenable),                               //                                          .byteenable
		.nios2_cpu_data_master_read                      (nios2_cpu_data_master_read),                                     //                                          .read
		.nios2_cpu_data_master_readdata                  (nios2_cpu_data_master_readdata),                                 //                                          .readdata
		.nios2_cpu_data_master_write                     (nios2_cpu_data_master_write),                                    //                                          .write
		.nios2_cpu_data_master_writedata                 (nios2_cpu_data_master_writedata),                                //                                          .writedata
		.nios2_cpu_data_master_debugaccess               (nios2_cpu_data_master_debugaccess),                              //                                          .debugaccess
		.nios2_cpu_instruction_master_address            (nios2_cpu_instruction_master_address),                           //              nios2_cpu_instruction_master.address
		.nios2_cpu_instruction_master_waitrequest        (nios2_cpu_instruction_master_waitrequest),                       //                                          .waitrequest
		.nios2_cpu_instruction_master_read               (nios2_cpu_instruction_master_read),                              //                                          .read
		.nios2_cpu_instruction_master_readdata           (nios2_cpu_instruction_master_readdata),                          //                                          .readdata
		.Av_FIFO_Int_0_avalon_slave_0_address            (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_address),         //              Av_FIFO_Int_0_avalon_slave_0.address
		.Av_FIFO_Int_0_avalon_slave_0_write              (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_write),           //                                          .write
		.Av_FIFO_Int_0_avalon_slave_0_read               (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_read),            //                                          .read
		.Av_FIFO_Int_0_avalon_slave_0_readdata           (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_readdata),        //                                          .readdata
		.Av_FIFO_Int_0_avalon_slave_0_writedata          (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_writedata),       //                                          .writedata
		.Av_FIFO_Int_0_avalon_slave_0_chipselect         (mm_interconnect_0_av_fifo_int_0_avalon_slave_0_chipselect),      //                                          .chipselect
		.dac_spi1_spi_control_port_address               (mm_interconnect_0_dac_spi1_spi_control_port_address),            //                 dac_spi1_spi_control_port.address
		.dac_spi1_spi_control_port_write                 (mm_interconnect_0_dac_spi1_spi_control_port_write),              //                                          .write
		.dac_spi1_spi_control_port_read                  (mm_interconnect_0_dac_spi1_spi_control_port_read),               //                                          .read
		.dac_spi1_spi_control_port_readdata              (mm_interconnect_0_dac_spi1_spi_control_port_readdata),           //                                          .readdata
		.dac_spi1_spi_control_port_writedata             (mm_interconnect_0_dac_spi1_spi_control_port_writedata),          //                                          .writedata
		.dac_spi1_spi_control_port_chipselect            (mm_interconnect_0_dac_spi1_spi_control_port_chipselect),         //                                          .chipselect
		.fpga_spi0_spi_control_port_address              (mm_interconnect_0_fpga_spi0_spi_control_port_address),           //                fpga_spi0_spi_control_port.address
		.fpga_spi0_spi_control_port_write                (mm_interconnect_0_fpga_spi0_spi_control_port_write),             //                                          .write
		.fpga_spi0_spi_control_port_read                 (mm_interconnect_0_fpga_spi0_spi_control_port_read),              //                                          .read
		.fpga_spi0_spi_control_port_readdata             (mm_interconnect_0_fpga_spi0_spi_control_port_readdata),          //                                          .readdata
		.fpga_spi0_spi_control_port_writedata            (mm_interconnect_0_fpga_spi0_spi_control_port_writedata),         //                                          .writedata
		.fpga_spi0_spi_control_port_chipselect           (mm_interconnect_0_fpga_spi0_spi_control_port_chipselect),        //                                          .chipselect
		.gpi_0_s1_address                                (mm_interconnect_0_gpi_0_s1_address),                             //                                  gpi_0_s1.address
		.gpi_0_s1_readdata                               (mm_interconnect_0_gpi_0_s1_readdata),                            //                                          .readdata
		.gpio_0_s1_address                               (mm_interconnect_0_gpio_0_s1_address),                            //                                 gpio_0_s1.address
		.gpio_0_s1_write                                 (mm_interconnect_0_gpio_0_s1_write),                              //                                          .write
		.gpio_0_s1_readdata                              (mm_interconnect_0_gpio_0_s1_readdata),                           //                                          .readdata
		.gpio_0_s1_writedata                             (mm_interconnect_0_gpio_0_s1_writedata),                          //                                          .writedata
		.gpio_0_s1_chipselect                            (mm_interconnect_0_gpio_0_s1_chipselect),                         //                                          .chipselect
		.i2c_opencores_0_avalon_slave_0_address          (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_address),       //            i2c_opencores_0_avalon_slave_0.address
		.i2c_opencores_0_avalon_slave_0_write            (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_write),         //                                          .write
		.i2c_opencores_0_avalon_slave_0_readdata         (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_readdata),      //                                          .readdata
		.i2c_opencores_0_avalon_slave_0_writedata        (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_writedata),     //                                          .writedata
		.i2c_opencores_0_avalon_slave_0_waitrequest      (~mm_interconnect_0_i2c_opencores_0_avalon_slave_0_waitrequest),  //                                          .waitrequest
		.i2c_opencores_0_avalon_slave_0_chipselect       (mm_interconnect_0_i2c_opencores_0_avalon_slave_0_chipselect),    //                                          .chipselect
		.jtag_uart_0_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),        //             jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),          //                                          .write
		.jtag_uart_0_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),           //                                          .read
		.jtag_uart_0_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),       //                                          .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),      //                                          .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),    //                                          .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),     //                                          .chipselect
		.nios2_cpu_debug_mem_slave_address               (mm_interconnect_0_nios2_cpu_debug_mem_slave_address),            //                 nios2_cpu_debug_mem_slave.address
		.nios2_cpu_debug_mem_slave_write                 (mm_interconnect_0_nios2_cpu_debug_mem_slave_write),              //                                          .write
		.nios2_cpu_debug_mem_slave_read                  (mm_interconnect_0_nios2_cpu_debug_mem_slave_read),               //                                          .read
		.nios2_cpu_debug_mem_slave_readdata              (mm_interconnect_0_nios2_cpu_debug_mem_slave_readdata),           //                                          .readdata
		.nios2_cpu_debug_mem_slave_writedata             (mm_interconnect_0_nios2_cpu_debug_mem_slave_writedata),          //                                          .writedata
		.nios2_cpu_debug_mem_slave_byteenable            (mm_interconnect_0_nios2_cpu_debug_mem_slave_byteenable),         //                                          .byteenable
		.nios2_cpu_debug_mem_slave_waitrequest           (mm_interconnect_0_nios2_cpu_debug_mem_slave_waitrequest),        //                                          .waitrequest
		.nios2_cpu_debug_mem_slave_debugaccess           (mm_interconnect_0_nios2_cpu_debug_mem_slave_debugaccess),        //                                          .debugaccess
		.oc_mem_s1_address                               (mm_interconnect_0_oc_mem_s1_address),                            //                                 oc_mem_s1.address
		.oc_mem_s1_write                                 (mm_interconnect_0_oc_mem_s1_write),                              //                                          .write
		.oc_mem_s1_readdata                              (mm_interconnect_0_oc_mem_s1_readdata),                           //                                          .readdata
		.oc_mem_s1_writedata                             (mm_interconnect_0_oc_mem_s1_writedata),                          //                                          .writedata
		.oc_mem_s1_byteenable                            (mm_interconnect_0_oc_mem_s1_byteenable),                         //                                          .byteenable
		.oc_mem_s1_chipselect                            (mm_interconnect_0_oc_mem_s1_chipselect),                         //                                          .chipselect
		.oc_mem_s1_clken                                 (mm_interconnect_0_oc_mem_s1_clken),                              //                                          .clken
		.pll_reconfig_0_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_address),     //          pll_reconfig_0_mgmt_avalon_slave.address
		.pll_reconfig_0_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_0_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_0_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_0_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_0_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_0_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.pll_reconfig_1_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_address),     //          pll_reconfig_1_mgmt_avalon_slave.address
		.pll_reconfig_1_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_1_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_1_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_1_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_1_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_1_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.pll_reconfig_2_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_address),     //          pll_reconfig_2_mgmt_avalon_slave.address
		.pll_reconfig_2_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_2_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_2_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_2_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_2_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_2_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.pll_reconfig_3_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_address),     //          pll_reconfig_3_mgmt_avalon_slave.address
		.pll_reconfig_3_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_3_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_3_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_3_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_3_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_3_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.pll_reconfig_4_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_address),     //          pll_reconfig_4_mgmt_avalon_slave.address
		.pll_reconfig_4_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_4_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_4_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_4_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_4_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_4_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.pll_reconfig_5_mgmt_avalon_slave_address        (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_address),     //          pll_reconfig_5_mgmt_avalon_slave.address
		.pll_reconfig_5_mgmt_avalon_slave_write          (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_write),       //                                          .write
		.pll_reconfig_5_mgmt_avalon_slave_read           (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_read),        //                                          .read
		.pll_reconfig_5_mgmt_avalon_slave_readdata       (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_readdata),    //                                          .readdata
		.pll_reconfig_5_mgmt_avalon_slave_writedata      (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_writedata),   //                                          .writedata
		.pll_reconfig_5_mgmt_avalon_slave_waitrequest    (mm_interconnect_0_pll_reconfig_5_mgmt_avalon_slave_waitrequest), //                                          .waitrequest
		.PLL_RST_s1_address                              (mm_interconnect_0_pll_rst_s1_address),                           //                                PLL_RST_s1.address
		.PLL_RST_s1_write                                (mm_interconnect_0_pll_rst_s1_write),                             //                                          .write
		.PLL_RST_s1_readdata                             (mm_interconnect_0_pll_rst_s1_readdata),                          //                                          .readdata
		.PLL_RST_s1_writedata                            (mm_interconnect_0_pll_rst_s1_writedata),                         //                                          .writedata
		.PLL_RST_s1_chipselect                           (mm_interconnect_0_pll_rst_s1_chipselect),                        //                                          .chipselect
		.PLLCFG_Command_s1_address                       (mm_interconnect_0_pllcfg_command_s1_address),                    //                         PLLCFG_Command_s1.address
		.PLLCFG_Command_s1_readdata                      (mm_interconnect_0_pllcfg_command_s1_readdata),                   //                                          .readdata
		.PLLCFG_SPI_spi_control_port_address             (mm_interconnect_0_pllcfg_spi_spi_control_port_address),          //               PLLCFG_SPI_spi_control_port.address
		.PLLCFG_SPI_spi_control_port_write               (mm_interconnect_0_pllcfg_spi_spi_control_port_write),            //                                          .write
		.PLLCFG_SPI_spi_control_port_read                (mm_interconnect_0_pllcfg_spi_spi_control_port_read),             //                                          .read
		.PLLCFG_SPI_spi_control_port_readdata            (mm_interconnect_0_pllcfg_spi_spi_control_port_readdata),         //                                          .readdata
		.PLLCFG_SPI_spi_control_port_writedata           (mm_interconnect_0_pllcfg_spi_spi_control_port_writedata),        //                                          .writedata
		.PLLCFG_SPI_spi_control_port_chipselect          (mm_interconnect_0_pllcfg_spi_spi_control_port_chipselect),       //                                          .chipselect
		.PLLCFG_Status_s1_address                        (mm_interconnect_0_pllcfg_status_s1_address),                     //                          PLLCFG_Status_s1.address
		.PLLCFG_Status_s1_write                          (mm_interconnect_0_pllcfg_status_s1_write),                       //                                          .write
		.PLLCFG_Status_s1_readdata                       (mm_interconnect_0_pllcfg_status_s1_readdata),                    //                                          .readdata
		.PLLCFG_Status_s1_writedata                      (mm_interconnect_0_pllcfg_status_s1_writedata),                   //                                          .writedata
		.PLLCFG_Status_s1_chipselect                     (mm_interconnect_0_pllcfg_status_s1_chipselect),                  //                                          .chipselect
		.sysid_qsys_0_control_slave_address              (mm_interconnect_0_sysid_qsys_0_control_slave_address),           //                sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata             (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)           //                                          .readdata
	);

	nios_cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_cpu_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_cpu_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_cpu_debug_reset_request_reset),    // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
