-- ddr3_av_x64_tester.vhd

-- Generated using ACDS version 16.1 200

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ddr3_av_x64_tester is
	port (
		avl_ready           : in  std_logic                     := '0';             --       avl.waitrequest_n
		avl_addr            : out std_logic_vector(25 downto 0);                    --          .address
		avl_size            : out std_logic_vector(1 downto 0);                     --          .burstcount
		avl_wdata           : out std_logic_vector(63 downto 0);                    --          .writedata
		avl_rdata           : in  std_logic_vector(63 downto 0) := (others => '0'); --          .readdata
		avl_write_req       : out std_logic;                                        --          .write
		avl_read_req        : out std_logic;                                        --          .read
		avl_rdata_valid     : in  std_logic                     := '0';             --          .readdatavalid
		avl_be              : out std_logic_vector(7 downto 0);                     --          .byteenable
		avl_burstbegin      : out std_logic;                                        --          .beginbursttransfer
		clk                 : in  std_logic                     := '0';             -- avl_clock.clk
		reset_n             : in  std_logic                     := '0';             -- avl_reset.reset_n
		pnf_per_bit         : out std_logic_vector(63 downto 0);                    --       pnf.pnf_per_bit
		pnf_per_bit_persist : out std_logic_vector(63 downto 0);                    --          .pnf_per_bit_persist
		pass                : out std_logic;                                        --    status.pass
		fail                : out std_logic;                                        --          .fail
		test_complete       : out std_logic                                         --          .test_complete
	);
end entity ddr3_av_x64_tester;

architecture rtl of ddr3_av_x64_tester is
	component ddr3_av_x64_tester_mm_traffic_generator_0 is
		generic (
			DEVICE_FAMILY                          : string  := "";
			TG_AVL_DATA_WIDTH                      : integer := 32;
			TG_AVL_ADDR_WIDTH                      : integer := 25;
			TG_AVL_WORD_ADDR_WIDTH                 : integer := 25;
			TG_AVL_SIZE_WIDTH                      : integer := 2;
			TG_AVL_BE_WIDTH                        : integer := 2;
			DRIVER_SIGNATURE                       : integer := 0;
			TG_GEN_BYTE_ADDR                       : boolean := true;
			TG_NUM_DRIVER_LOOP                     : integer := 1000;
			TG_ENABLE_UNIX_ID                      : boolean := false;
			TG_USE_UNIX_ID                         : integer := 0;
			TG_RANDOM_BYTE_ENABLE                  : boolean := false;
			TG_ENABLE_READ_COMPARE                 : boolean := true;
			TG_POWER_OF_TWO_BURSTS_ONLY            : boolean := false;
			TG_BURST_ON_BURST_BOUNDARY             : boolean := false;
			TG_DO_NOT_CROSS_4KB_BOUNDARY           : boolean := false;
			TG_TIMEOUT_COUNTER_WIDTH               : integer := 32;
			TG_MAX_READ_LATENCY                    : integer := 20;
			TG_SINGLE_RW_SEQ_ADDR_COUNT            : integer := 32;
			TG_SINGLE_RW_RAND_ADDR_COUNT           : integer := 32;
			TG_SINGLE_RW_RAND_SEQ_ADDR_COUNT       : integer := 32;
			TG_BLOCK_RW_SEQ_ADDR_COUNT             : integer := 8;
			TG_BLOCK_RW_RAND_ADDR_COUNT            : integer := 8;
			TG_BLOCK_RW_RAND_SEQ_ADDR_COUNT        : integer := 8;
			TG_BLOCK_RW_BLOCK_SIZE                 : integer := 8;
			TG_TEMPLATE_STAGE_COUNT                : integer := 4;
			TG_SEQ_ADDR_GEN_MIN_BURSTCOUNT         : integer := 1;
			TG_SEQ_ADDR_GEN_MAX_BURSTCOUNT         : integer := 2;
			TG_RAND_ADDR_GEN_MIN_BURSTCOUNT        : integer := 1;
			TG_RAND_ADDR_GEN_MAX_BURSTCOUNT        : integer := 2;
			TG_RAND_SEQ_ADDR_GEN_MIN_BURSTCOUNT    : integer := 1;
			TG_RAND_SEQ_ADDR_GEN_MAX_BURSTCOUNT    : integer := 2;
			TG_RAND_SEQ_ADDR_GEN_RAND_ADDR_PERCENT : integer := 50
		);
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset_n             : in  std_logic                     := 'X';             -- reset_n
			pass                : out std_logic;                                        -- pass
			fail                : out std_logic;                                        -- fail
			test_complete       : out std_logic;                                        -- test_complete
			pnf_per_bit         : out std_logic_vector(63 downto 0);                    -- pnf_per_bit
			pnf_per_bit_persist : out std_logic_vector(63 downto 0);                    -- pnf_per_bit_persist
			avl_ready           : in  std_logic                     := 'X';             -- waitrequest_n
			avl_addr            : out std_logic_vector(25 downto 0);                    -- address
			avl_size            : out std_logic_vector(1 downto 0);                     -- burstcount
			avl_wdata           : out std_logic_vector(63 downto 0);                    -- writedata
			avl_rdata           : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			avl_write_req       : out std_logic;                                        -- write
			avl_read_req        : out std_logic;                                        -- read
			avl_rdata_valid     : in  std_logic                     := 'X';             -- readdatavalid
			avl_be              : out std_logic_vector(7 downto 0);                     -- byteenable
			avl_burstbegin      : out std_logic                                         -- beginbursttransfer
		);
	end component ddr3_av_x64_tester_mm_traffic_generator_0;

begin

	mm_traffic_generator_0 : component ddr3_av_x64_tester_mm_traffic_generator_0
		generic map (
			DEVICE_FAMILY                          => "Cyclone V",
			TG_AVL_DATA_WIDTH                      => 64,
			TG_AVL_ADDR_WIDTH                      => 26,
			TG_AVL_WORD_ADDR_WIDTH                 => 23,
			TG_AVL_SIZE_WIDTH                      => 2,
			TG_AVL_BE_WIDTH                        => 8,
			DRIVER_SIGNATURE                       => 1431634081,
			TG_GEN_BYTE_ADDR                       => true,
			TG_NUM_DRIVER_LOOP                     => 1000,
			TG_ENABLE_UNIX_ID                      => false,
			TG_USE_UNIX_ID                         => 0,
			TG_RANDOM_BYTE_ENABLE                  => false,
			TG_ENABLE_READ_COMPARE                 => true,
			TG_POWER_OF_TWO_BURSTS_ONLY            => false,
			TG_BURST_ON_BURST_BOUNDARY             => false,
			TG_DO_NOT_CROSS_4KB_BOUNDARY           => false,
			TG_TIMEOUT_COUNTER_WIDTH               => 32,
			TG_MAX_READ_LATENCY                    => 20,
			TG_SINGLE_RW_SEQ_ADDR_COUNT            => 32,
			TG_SINGLE_RW_RAND_ADDR_COUNT           => 32,
			TG_SINGLE_RW_RAND_SEQ_ADDR_COUNT       => 32,
			TG_BLOCK_RW_SEQ_ADDR_COUNT             => 8,
			TG_BLOCK_RW_RAND_ADDR_COUNT            => 8,
			TG_BLOCK_RW_RAND_SEQ_ADDR_COUNT        => 8,
			TG_BLOCK_RW_BLOCK_SIZE                 => 8,
			TG_TEMPLATE_STAGE_COUNT                => 4,
			TG_SEQ_ADDR_GEN_MIN_BURSTCOUNT         => 1,
			TG_SEQ_ADDR_GEN_MAX_BURSTCOUNT         => 2,
			TG_RAND_ADDR_GEN_MIN_BURSTCOUNT        => 1,
			TG_RAND_ADDR_GEN_MAX_BURSTCOUNT        => 2,
			TG_RAND_SEQ_ADDR_GEN_MIN_BURSTCOUNT    => 1,
			TG_RAND_SEQ_ADDR_GEN_MAX_BURSTCOUNT    => 2,
			TG_RAND_SEQ_ADDR_GEN_RAND_ADDR_PERCENT => 50
		)
		port map (
			clk                 => clk,                 -- avl_clock.clk
			reset_n             => reset_n,             -- avl_reset.reset_n
			pass                => pass,                --    status.pass
			fail                => fail,                --          .fail
			test_complete       => test_complete,       --          .test_complete
			pnf_per_bit         => pnf_per_bit,         --       pnf.pnf_per_bit
			pnf_per_bit_persist => pnf_per_bit_persist, --          .pnf_per_bit_persist
			avl_ready           => avl_ready,           --       avl.waitrequest_n
			avl_addr            => avl_addr,            --          .address
			avl_size            => avl_size,            --          .burstcount
			avl_wdata           => avl_wdata,           --          .writedata
			avl_rdata           => avl_rdata,           --          .readdata
			avl_write_req       => avl_write_req,       --          .write
			avl_read_req        => avl_read_req,        --          .read
			avl_rdata_valid     => avl_rdata_valid,     --          .readdatavalid
			avl_be              => avl_be,              --          .byteenable
			avl_burstbegin      => avl_burstbegin       --          .beginbursttransfer
		);

end architecture rtl; -- of ddr3_av_x64_tester
